`define R_ins 7'b0110011

`define J_ins 7'b1101111
`define B_ins 7'b1100011
`define S_ins 7'b0100011

`define I_ins_J 7'b1100111
`define I_ins_R 7'b0010011
`define I_ins_L 7'b0000011

`define U_ins_lui   7'b0110111
`define U_ins_auipc 7'b0010111

`define ADD 	4'b0000
`define SUB 	4'b0001
`define SLL 	4'b0010
`define SLT 	4'b0011
`define SLTU	4'b0100
`define SRA 	4'b0101
`define OR 	    4'b0111
`define AND 	4'b1000
`define XOR 	4'b1001
`define SRL     4'b1011 

`define SB      3'b000 
`define SH      3'b001 
`define SW      3'b010 

`define BEQ     3'b000
`define BNE     3'b001
`define BLT     3'b010
`define BGE     3'b011
`define BLTU    3'b100
`define BGEU    3'b101


   
`define COMPARE 4'b1111   
                  
                  
                  
                  
                  
